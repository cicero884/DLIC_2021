module traffic_light (
  input  clk,
  input  rst,
  input  pass,
  output R,
  output G,
  output Y
);

endmodule
